//--------------------------------------
//-- SinTable.vhd
//-- Written by Gadi and Eran Tuchman.
//-- All rights reserved, Copyright 2009
//-- SystemVerilog version June 2018 Alex Grinshpun
//--------------------------------------


module	sintable	 #(
					COUNT_SIZE = 8
		)	
		(	
//		--////////////////////	Clock Input	 	////////////////////	
					input		logic	CLK,
					input		logic	RESETn,
					input		logic [COUNT_SIZE-1:0]	ADDR,
					output	logic [15:0]	Q
			);






localparam int table_size = (2**COUNT_SIZE)-1;


const logic [0:table_size-1] [15:0] sin_table = {

16'h0000,
16'h0188,
16'h0311,
16'h0499,
16'h0620,
16'h07A6,
16'h092B,
16'h0AAF,
16'h0C31,
16'h0DB1,
16'h0F2F,
16'h10AB,
16'h1224,
16'h139A,
16'h150E,
16'h167E,
16'h17EA,
16'h1953,
16'h1AB8,
16'h1C19,
16'h1D76,
16'h1ECE,
16'h2021,
16'h216F,
16'h22B9,
16'h23FC,
16'h253B,
16'h2673,
16'h27A6,
16'h28D2,
16'h29F8,
16'h2B18,
16'h2C31,
16'h2D43,
16'h2E4F,
16'h2F53,
16'h3050,
16'h3145,
16'h3233,
16'h3319,
16'h33F7,
16'h34CD,
16'h359B,
16'h3661,
16'h371E,
16'h37D3,
16'h387F,
16'h3923,
16'h39BE,
16'h3A4F,
16'h3AD8,
16'h3B58,
16'h3BCF,
16'h3C3C,
16'h3CA0,
16'h3CFB,
16'h3D4C,
16'h3D94,
16'h3DD2,
16'h3E07,
16'h3E32,
16'h3E54,
16'h3E6C,
16'h3E7B,
16'h3E80,
16'h3E7B,
16'h3E6C,
16'h3E54,
16'h3E32,
16'h3E07,
16'h3DD2,
16'h3D94,
16'h3D4C,
16'h3CFB,
16'h3CA0,
16'h3C3C,
16'h3BCF,
16'h3B58,
16'h3AD8,
16'h3A4F,
16'h39BE,
16'h3923,
16'h387F,
16'h37D3,
16'h371E,
16'h3661,
16'h359B,
16'h34CD,
16'h33F7,
16'h3319,
16'h3233,
16'h3145,
16'h3050,
16'h2F53,
16'h2E4F,
16'h2D43,
16'h2C31,
16'h2B18,
16'h29F8,
16'h28D2,
16'h27A6,
16'h2673,
16'h253B,
16'h23FC,
16'h22B9,
16'h216F,
16'h2021,
16'h1ECE,
16'h1D76,
16'h1C19,
16'h1AB8,
16'h1953,
16'h17EA,
16'h167E,
16'h150E,
16'h139A,
16'h1224,
16'h10AB,
16'h0F2F,
16'h0DB1,
16'h0C31,
16'h0AAF,
16'h092B,
16'h07A6,
16'h0620,
16'h0499,
16'h0311,
16'h0188,
16'h0000,
16'hFE78,
16'hFCEF,
16'hFB67,
16'hF9E0,
16'hF85A,
16'hF6D5,
16'hF551,
16'hF3CF,
16'hF24F,
16'hF0D1,
16'hEF55,
16'hEDDC,
16'hEC66,
16'hEAF2,
16'hE982,
16'hE816,
16'hE6AD,
16'hE548,
16'hE3E7,
16'hE28A,
16'hE132,
16'hDFDF,
16'hDE91,
16'hDD47,
16'hDC04,
16'hDAC5,
16'hD98D,
16'hD85A,
16'hD72E,
16'hD608,
16'hD4E8,
16'hD3CF,
16'hD2BD,
16'hD1B1,
16'hD0AD,
16'hCFB0,
16'hCEBB,
16'hCDCD,
16'hCCE7,
16'hCC09,
16'hCB33,
16'hCA65,
16'hC99F,
16'hC8E2,
16'hC82D,
16'hC781,
16'hC6DD,
16'hC642,
16'hC5B1,
16'hC528,
16'hC4A8,
16'hC431,
16'hC3C4,
16'hC360,
16'hC305,
16'hC2B4,
16'hC26C,
16'hC22E,
16'hC1F9,
16'hC1CE,
16'hC1AC,
16'hC194,
16'hC185,
16'hC180,
16'hC185,
16'hC194,
16'hC1AC,
16'hC1CE,
16'hC1F9,
16'hC22E,
16'hC26C,
16'hC2B4,
16'hC305,
16'hC360,
16'hC3C4,
16'hC431,
16'hC4A8,
16'hC528,
16'hC5B1,
16'hC642,
16'hC6DD,
16'hC781,
16'hC82D,
16'hC8E2,
16'hC99F,
16'hCA65,
16'hCB33,
16'hCC09,
16'hCCE7,
16'hCDCD,
16'hCEBB,
16'hCFB0,
16'hD0AD,
16'hD1B1,
16'hD2BD,
16'hD3CF,
16'hD4E8,
16'hD608,
16'hD72E,
16'hD85A,
16'hD98D,
16'hDAC5,
16'hDC04,
16'hDD47,
16'hDE91,
16'hDFDF,
16'hE132,
16'hE28A,
16'hE3E7,
16'hE548,
16'hE6AD,
16'hE816,
16'hE982,
16'hEAF2,
16'hEC66,
16'hEDDC,
16'hEF55,
16'hF0D1,
16'hF24F,
16'hF3CF,
16'hF551,
16'hF6D5,
16'hF85A,
16'hF9E0,
16'hFB67,
16'hFCEF,
16'hFE78
 };

 

always_ff@(posedge CLK or negedge RESETn)
begin
	if(!RESETn)
	begin
		Q	<= 16'h0;
	end
	else 
		Q	<= sin_table[ADDR];

end
endmodule
